module not_gate_st ( input a , output y) ;
	assign y=not(a,y); 
endmodule