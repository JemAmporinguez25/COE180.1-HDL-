
module not_gate_df(input a,output y); // define module to test run
	assign y=~a ;
endmodule
