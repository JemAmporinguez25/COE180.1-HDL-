module and_gate_st ( input a , b , output y) ;
	and(a , b , y );
endmodule