module or_gate_st ( input a , b , output y) ;
	or(y , a , b );
	
endmodule